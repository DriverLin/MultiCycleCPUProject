//////////////////////////////////////////////////////////////////////////////////
// 模块名称: IM
// 模块功能: 指令存储器
//          存储指令
//////////////////////////////////////////////////////////////////////////////////
module IM(
    input               clk,
    input	[11:2]      addr,
    output	reg[31:0]   dout
);
    reg     [31:0]  ROM[1023:0];
    initial begin
ROM[0] = 0'b00000001010010100100100000100010;
ROM[1] = 0'b00100001001010010000000000000001;
ROM[2] = 0'b00001000000000000000000000000001;
    end
    always @(posedge clk) begin
        dout = ROM[addr[11:2]][31:0];
    end
endmodule
